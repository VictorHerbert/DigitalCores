/*package vga_config;

    typedef struct {
        int red;
        int green;
        int blue;
        
        int width;
    } PixelWidth;

    typedef struct {
        int visible_area;
        int front_porch;
        int sync_pulse;
        int back_porch;

        int line;
    } VGADimentionTiming;

    typedef struct {
        VGADimentionTiming horizontal;
        VGADimentionTiming vertical;
        int mem_size;
    } VGATiming;

endpackage*/



